module tb_uart_top;

  logic pclk = 0;
  logic presetn;
  logic psel;
  logic penable;
  logic pwrite;
  logic [31:0] paddr;
  logic [31:0] pwdata;
  
  logic uart_rxd;
  
  logic pready;
  logic [31:0] prdata;
  
  logic uart_txd;

  always #5 pclk = ~ pclk;

  uart_top u_uart_top (
   .pclk       ( pclk       ),
   .presetn    ( presetn    ),
   .psel       ( psel       ),
   .penable    ( penable    ),
   .pwrite     ( pwrite     ),
   .paddr      ( paddr      ),
   .pwdata     ( pwdata     ),
   
   .uart_rxd   ( uart_rxd   ),
   
   .pready     ( pready     ),
   .prdata     ( prdata     ),
   
   .uart_txd    ( uart_txd    ),
   .uart_intpt ( uart_intpt )
  );


  //..............reset...................
  task reset;
    presetn = 1'b0;
    @(posedge pclk);
    presetn = 1'b1;
  endtask
  //......................................


  initial begin

    presetn  = 0;
    psel     = 0;
    penable  = 0;
    pwrite   = 0;
    paddr    = 32'h0;
    pwdata   = 32'h0;
    uart_rxd = 0;
    repeat(4) @(posedge pclk);
    reset;

    repeat(40) @(posedge pclk);

    dll_wr(8'b011);
    write(32'h8,{24'b0,8'b00000001}); // FCR -> fifen = 1
    
    lcr_wr(8'b10111111);
    //write(32'h8,{24'b0,8'b00000001}); // FCR -> fifen = 1
    thr_wr(8'b11110011);
    thr_wr(8'b11111111);
    thr_wr(8'b00001000);
    thr_wr(8'b10000001);
    thr_wr(8'b00000000);
    
    
    pwm (1,1);     
    
    

    #200000;


    $finish;
  end
  
  task thr_wr (input [7:0] transmit_data);
    begin 
      @(posedge pclk);
      psel = 1;
      pwrite = 1;
      paddr = 32'h0;
      pwdata = {24'b0,transmit_data};
      @(posedge pclk);  
      penable = 1;   
      @(posedge pclk);
      psel = 0;
      pwrite = 0;
      penable = 0; 
    end
  endtask  

  task dll_wr (input [7:0] divisor_l);
    begin 
      @(posedge pclk);
      psel = 1;
      pwrite = 1;
      paddr = 32'h0020;
      pwdata = {24'b0,divisor_l};
      @(posedge pclk);  
      penable = 1;   
      @(posedge pclk);
      psel = 0;
      pwrite = 0;
      penable = 0; 
    end
  endtask

  task lcr_wr (input [7:0] line_control);
    begin 
      @(posedge pclk);
      psel = 1;
      pwrite = 1;
      paddr = 32'h000C;
      pwdata = {24'b0,line_control};
      @(posedge pclk);  
      penable = 1;   
      @(posedge pclk);
      psel = 0;
      pwrite = 0;
      penable = 0; 
    end
  endtask
  
  task write (input [31:0] adr, input [31:0] data );
    begin 
      @(posedge pclk);
      psel = 1;
      pwrite = 1;
      paddr = adr;
      pwdata = data;
      @(posedge pclk);  
      penable = 1;   
      @(posedge pclk);
      psel = 0;
      pwrite = 0;
      penable = 0; 
    end
  endtask

  task pwm (input tx_en, input rx_en);
    begin 
      @(posedge pclk);
      psel = 1;
      pwrite = 1;
      paddr = 32'h0030;
      pwdata = {32'hFFFFFFFF};
      @(posedge pclk);  
      penable = 1;   
      @(posedge pclk);
      psel = 0;
      pwrite = 0;
      penable = 0; 
    end
  endtask

endmodule